package My_Package;
import uvm_pkg::*;
`include "uvm_macros.svh"

`include "My_Sequence_Item.sv"
`include "My_Sequence.sv"
`include "My_Driver.sv"
`include "My_Monitor.sv"
`include "My_Sequencer.sv"
`include "My_Agent.sv"
`include "My_Scoreboard.sv"
`include "My_Subscriber.sv"
`include "My_Environment.sv"
`include "My_Test.sv"

endpackage : My_Package